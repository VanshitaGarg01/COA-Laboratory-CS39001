module branch_unit (
    input nextPC,
    
);
    
endmodule
