module datapath (
    
);
    
endmodule