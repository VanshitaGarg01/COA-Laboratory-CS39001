module instruction_memory (pc, instruction, clk, rst);
    input clk, rst;
    input [31:0] pc;
    output [31:0] instruction;
    // instruction_memory instantiate
endmodule