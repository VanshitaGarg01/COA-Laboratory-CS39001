module pc (
    input next_inst_addr,
    input clk, 
    input rst,
    output inst_addr
);

    always @(posedge clk or posedge rst) begin
        
    end

endmodule
